library verilog;
use verilog.vl_types.all;
entity TB_regis is
end TB_regis;
