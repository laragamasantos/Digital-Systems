library verilog;
use verilog.vl_types.all;
entity contador_4bits_tb is
end contador_4bits_tb;
