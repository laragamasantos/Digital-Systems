library verilog;
use verilog.vl_types.all;
entity exemplo_ou is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        S               : out    vl_logic
    );
end exemplo_ou;
