library verilog;
use verilog.vl_types.all;
entity contador_sincrono_tb is
end contador_sincrono_tb;
